module cputop(
    input clk,
    input rst_n,
    output [31:0] instrmem_instr_addr,
    input [31:0] instrmem_instr_data,
    output datamem_r_en,
    input [31:0] datamem_datar,
    output datamem_w_en,
    output [31:0] datamem_dataw
)；
endmodule